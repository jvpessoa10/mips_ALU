module mux(i)