module ALUControl(
	input [5:0] funct,
	input [1:0] ALUOp,
	output [3:0] Operation
);


endmodule